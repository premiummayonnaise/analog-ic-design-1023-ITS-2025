** sch_path: /foss/designs/analog-ic-design-1023-ITS-2025/week01_mosfet_cmos/tugas1_iv_curve/mosfet-iv-characteristics.sch
**.subckt mosfet-iv-characteristics
V1 VGS GND 0
V2 VDS GND 3.3
XM1 VDS VGS GND GND nfet_03v3_dss L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
**** begin user architecture code

.include /foss/pdks/gf180mcuD/libs.tech/ngspice/design.ngspice
.lib /foss/pdks/gf180mcuD/libs.tech/ngspice/sm141064.ngspice typical
.lib /foss/pdks/gf180mcuD/libs.tech/ngspice/smbb000149.ngspice typical




.control

	dc V2 0 3.3 0.01 V1 0 3.3 0.3
	plot -i(V2)

save all


.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
